module pipeline_reg #(
    parameter int DATA_WIDTH = 32
) (
    input  logic                   clk,
    input  logic                   rst_n,
    input  logic                   in_valid,
    output logic                   in_ready,
    input  logic [DATA_WIDTH-1:0]  in_data,
    output logic                   out_valid,
    input  logic                   out_ready,
    output logic [DATA_WIDTH-1:0]  out_data
);

    logic full;
    logic [DATA_WIDTH-1:0]  data_reg;
  
    assign in_ready  = ~full || out_ready;
    assign out_valid = full;
    assign out_data  = data_reg;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            full     <= 1'b0;
            data_reg <= '0;
        end
        else begin
          
            if (in_valid && in_ready) begin
                data_reg <= in_data;
                full     <= 1'b1;
            end
   
            else if (out_ready && full) begin
                full <= 1'b0;
            end
        end
    end

endmodule
